module
not_gate (
    input wire a,      // Input signal a
    output wire out    // Output signal
);

    // NOT gate logic
    assign out = ~a;

endmodule
